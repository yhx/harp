module array_accu_pl #(CACHE_WIDTH = 512, DATA_WIDTH = 32)
	(
		input clk,
		input rst,
		input inc,
		input [CACHE_WIDTH-1:0] array,
		output [CACHE_WIDTH-1:0] res,
		output ready
	);

	localparam DATA_SIZE = CACHE_WIDTH/DATA_WIDTH;

	reg [CACHE_WIDTH-1:0] add_0_res;

	assign res = add_0_res;

	reg enable0;
	assign ready = enable0 && !inc;

	always@(posedge clk)
	begin
		enable0 <= rst ? 1'b0 : inc;
	end

	genvar i;
	generate for (i=0; i<DATA_SIZE; i++)
		begin:adder
			always@(posedge clk)
			begin
				if (rst)
				begin
					add_0_res <= 0;
				end
				else if (inc)
				begin
					add_0_res[i<<5 +: DATA_WIDTH] <= array[i<<5 +: DATA_WIDTH] + add_0_res[i<<5 +: DATA_WIDTH];
				end
				else
				begin
					//$display("ADD_RES: %d@%d, %d@%d", add_3_res[0], 0, add_3_res[1], 1);
					add_0_res[i<<5 +: DATA_WIDTH] <= array[i<<5 +: DATA_WIDTH];
				end
			end
		end
	endgenerate

endmodule

