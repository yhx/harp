module conv2d
	(
		input [511:0] data;
		input [511:0] kernel;

		output [31:0] res;
	);


reg [511:0] buffer;

endmodule
